magic
tech scmos
timestamp 1710979321
<< ntransistor >>
rect 4 -1 6 3
rect 26 -1 28 3
rect 44 -1 46 3
<< ptransistor >>
rect 4 20 6 24
rect 26 20 28 24
rect 44 20 46 24
<< ndiffusion >>
rect 2 -1 4 3
rect 6 -1 14 3
rect 18 -1 26 3
rect 28 -1 30 3
rect 42 -1 44 3
rect 46 -1 47 3
<< pdiffusion >>
rect 2 20 4 24
rect 6 20 26 24
rect 28 20 30 24
rect 42 20 44 24
rect 46 20 47 24
<< ndcontact >>
rect -2 -1 2 3
rect 14 -1 18 3
rect 30 -1 34 3
rect 38 -1 42 3
rect 47 -1 51 3
<< pdcontact >>
rect -2 20 2 24
rect 30 20 34 24
rect 38 20 42 24
rect 47 20 51 24
<< psubstratepcontact >>
rect -2 -9 2 -5
rect 30 -9 34 -5
rect 38 -9 42 -5
<< nsubstratencontact >>
rect -2 28 2 32
rect 38 28 42 32
<< polysilicon >>
rect 4 24 6 26
rect 26 24 28 26
rect 44 24 46 26
rect 4 11 6 20
rect 26 19 28 20
rect 24 15 28 19
rect 2 7 6 11
rect 4 3 6 7
rect 26 3 28 15
rect 44 11 46 20
rect 42 7 46 11
rect 44 3 46 7
rect 4 -4 6 -1
rect 26 -3 28 -1
rect 44 -3 46 -1
<< polycontact >>
rect 20 15 24 19
rect -2 7 2 11
rect 38 7 42 11
<< metal1 >>
rect -4 28 -2 32
rect 2 28 38 32
rect 42 28 53 32
rect -2 24 2 28
rect 38 24 42 28
rect 30 11 34 20
rect 14 7 38 11
rect 14 3 18 7
rect 47 3 51 20
rect -2 -5 2 -1
rect 30 -5 34 -1
rect 38 -5 42 -1
rect -4 -9 -2 -5
rect 2 -9 30 -5
rect 34 -9 38 -5
rect 42 -9 54 -5
<< labels >>
rlabel polycontact 0 9 0 9 1 A
rlabel polycontact 40 9 40 9 1 INV
rlabel metal1 49 10 49 10 1 Y
rlabel psubstratepcontact 0 -7 0 -7 1 VSS
rlabel psubstratepcontact 32 -7 32 -7 1 VSS
rlabel psubstratepcontact 40 -7 40 -7 1 VSS
rlabel nsubstratencontact 0 30 0 30 1 VDD
rlabel nsubstratencontact 40 30 40 30 1 VDD
rlabel polycontact 22 17 22 17 1 B
<< end >>
