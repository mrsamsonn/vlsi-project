magic
tech scmos
timestamp 1709331696
<< ntransistor >>
rect 5 8 7 12
rect 16 8 18 12
rect 27 8 29 12
rect 38 8 40 12
rect 57 8 59 12
<< ptransistor >>
rect 5 41 7 45
rect 16 41 18 45
rect 27 41 29 45
rect 38 41 40 45
rect 57 41 59 45
<< ndiffusion >>
rect 4 8 5 12
rect 7 8 8 12
rect 12 8 16 12
rect 18 8 20 12
rect 24 8 27 12
rect 29 8 32 12
rect 36 8 38 12
rect 40 8 44 12
rect 56 8 57 12
rect 59 8 60 12
<< pdiffusion >>
rect 4 41 5 45
rect 7 41 16 45
rect 18 41 27 45
rect 29 41 38 45
rect 40 41 44 45
rect 56 41 57 45
rect 59 41 60 45
<< ndcontact >>
rect 0 8 4 12
rect 8 8 12 12
rect 20 8 24 12
rect 32 8 36 12
rect 44 8 48 12
rect 52 8 56 12
rect 60 8 64 12
<< pdcontact >>
rect 0 41 4 45
rect 44 41 48 45
rect 52 41 56 45
rect 60 41 64 45
<< psubstratepcontact >>
rect 8 0 12 4
rect 32 0 36 4
rect 52 0 56 4
<< nsubstratencontact >>
rect 0 49 4 53
rect 52 49 56 53
<< polysilicon >>
rect 5 45 7 47
rect 16 45 18 47
rect 27 45 29 47
rect 38 45 40 47
rect 57 45 59 47
rect 5 28 7 41
rect 16 28 18 41
rect 27 28 29 41
rect 38 28 40 41
rect 57 28 59 41
rect 4 24 7 28
rect 15 24 18 28
rect 26 24 29 28
rect 37 24 40 28
rect 56 24 59 28
rect 5 12 7 24
rect 16 12 18 24
rect 27 12 29 24
rect 38 12 40 24
rect 57 12 59 24
rect 5 6 7 8
rect 16 6 18 8
rect 27 6 29 8
rect 38 6 40 8
rect 57 6 59 8
<< polycontact >>
rect 0 24 4 28
rect 11 24 15 28
rect 22 24 26 28
rect 33 24 37 28
rect 52 24 56 28
<< metal1 >>
rect -4 49 0 53
rect 4 49 52 53
rect 0 45 4 49
rect 52 45 56 49
rect 44 28 48 41
rect 44 24 52 28
rect 44 20 48 24
rect 0 16 48 20
rect 0 12 4 16
rect 20 12 24 16
rect 44 12 48 16
rect 60 12 64 41
rect 8 4 12 8
rect 32 4 36 8
rect 52 4 56 8
rect 0 0 8 4
rect 12 0 32 4
rect 36 0 52 4
<< labels >>
rlabel metal1 -2 51 -2 51 4 VDD
rlabel metal1 2 2 2 2 1 VSS
rlabel polycontact 2 26 2 26 1 A
rlabel polycontact 13 26 13 26 1 B
rlabel polycontact 24 26 24 26 1 C
rlabel polycontact 35 26 35 26 1 D
rlabel polycontact 54 26 54 26 1 INV
rlabel metal1 62 26 62 26 7 Y
<< end >>
