magic
tech scmos
timestamp 1711427132
<< metal1 >>
rect 0 56 8 60
rect 266 28 272 32
rect 393 23 399 27
rect 0 0 8 4
rect 12 -8 16 -4
rect 185 -8 190 -4
rect 63 -25 67 -21
rect 152 -25 227 -21
rect 336 -24 344 -20
rect 152 -29 156 -25
rect 98 -33 156 -29
rect 168 -38 366 -34
<< m2contact >>
rect 366 28 370 32
rect 344 20 348 24
rect 94 12 98 16
rect 164 12 168 16
rect 332 12 336 16
rect 116 -16 120 -12
rect 332 -24 336 -20
rect 344 -24 348 -20
rect 94 -33 98 -29
rect 164 -38 168 -34
rect 366 -38 370 -34
<< metal2 >>
rect 94 -29 98 12
rect 164 -34 168 12
rect 332 -20 336 12
rect 344 -20 348 20
rect 366 -34 370 28
use 2or  2or_0
timestamp 1711420332
transform 1 0 346 0 1 9
box -10 -9 54 51
use half  half_0
timestamp 1711424539
transform 1 0 22 0 1 0
box -22 -25 148 60
use half  half_1
timestamp 1711424539
transform 1 0 190 0 1 0
box -22 -25 148 60
<< labels >>
rlabel metal1 398 25 398 25 1 Cout
rlabel metal1 270 30 270 30 1 Result
rlabel metal1 187 -6 187 -6 1 Cin
rlabel metal1 14 -6 14 -6 1 A
rlabel metal1 66 -23 66 -23 1 B
rlabel metal1 1 2 1 2 1 VSS
rlabel metal1 2 58 2 58 1 VDD
<< end >>
