magic
tech scmos
timestamp 1711410620
<< ntransistor >>
rect 6 8 8 12
rect 20 8 22 12
rect 43 8 45 12
rect 64 8 66 12
<< ptransistor >>
rect 6 40 8 44
rect 20 40 22 44
rect 43 40 45 44
rect 64 40 66 44
<< ndiffusion >>
rect 4 8 6 12
rect 8 8 20 12
rect 22 8 34 12
rect 38 8 43 12
rect 45 8 64 12
rect 66 8 70 12
<< pdiffusion >>
rect 4 40 6 44
rect 8 40 12 44
rect 16 40 20 44
rect 22 40 26 44
rect 38 40 43 44
rect 45 40 54 44
rect 58 40 64 44
rect 66 40 70 44
<< ndcontact >>
rect 0 8 4 12
rect 34 8 38 12
rect 70 8 74 12
<< pdcontact >>
rect 0 40 4 44
rect 12 40 16 44
rect 26 40 30 44
rect 34 40 38 44
rect 54 40 58 44
rect 70 40 74 44
<< psubstratepcontact >>
rect 34 0 38 4
<< nsubstratencontact >>
rect 12 56 16 60
<< polysilicon >>
rect 6 44 8 46
rect 20 44 22 46
rect 43 44 45 46
rect 64 44 66 46
rect 6 12 8 40
rect 20 12 22 40
rect 43 12 45 40
rect 64 12 66 40
rect 6 6 8 8
rect 20 6 22 8
rect 43 6 45 8
rect 64 6 66 8
<< polycontact >>
rect 2 25 6 29
rect 16 25 20 29
rect 39 25 43 29
rect 60 25 64 29
<< metal1 >>
rect -18 56 -12 60
rect -2 56 12 60
rect 16 56 80 60
rect 12 44 16 56
rect 26 48 58 52
rect 26 44 30 48
rect 54 44 58 48
rect 0 36 4 40
rect 26 36 30 40
rect 0 32 30 36
rect 34 36 38 40
rect 70 36 74 40
rect 34 32 74 36
rect -4 25 2 29
rect 70 28 82 32
rect 70 20 74 28
rect 0 16 74 20
rect 0 12 4 16
rect 70 12 74 16
rect 34 4 38 8
rect -18 0 -12 4
rect -2 0 34 4
rect 38 0 78 4
rect -12 -8 56 -4
rect 16 -16 92 -12
rect 39 -25 80 -21
<< m2contact >>
rect 12 25 16 29
rect 35 25 39 29
rect 56 25 60 29
rect -16 21 -12 25
rect 80 21 84 25
rect 92 8 96 12
rect -16 -8 -12 -4
rect 56 -8 60 -4
rect 12 -16 16 -12
rect 92 -16 96 -12
rect 35 -25 39 -21
rect 80 -25 84 -21
<< metal2 >>
rect -16 -4 -12 21
rect 12 -12 16 25
rect 35 -21 39 25
rect 56 -4 60 25
rect 80 -21 84 21
rect 92 -12 96 8
use INV  INV_1
timestamp 1711404725
transform 1 0 -13 0 1 -1
box -5 1 11 61
use INV  INV_2
timestamp 1711404725
transform 1 0 83 0 1 -1
box -5 1 11 61
<< labels >>
rlabel nsubstratencontact 14 58 14 58 5 VDD
rlabel polycontact 4 27 4 27 3 A
rlabel polycontact 18 27 18 27 1 B
rlabel metal1 -17 58 -17 58 1 VDD
rlabel metal1 -17 2 -17 2 1 VSS
rlabel psubstratepcontact 36 2 36 2 1 VSS
rlabel polycontact 41 27 41 27 1 B
rlabel polycontact 62 27 62 27 1 A
rlabel metal1 80 30 80 30 1 Y
<< end >>
