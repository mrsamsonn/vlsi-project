magic
tech scmos
timestamp 1711062510
<< ntransistor >>
rect 10 8 12 12
rect 20 8 22 12
<< ptransistor >>
rect 10 32 12 36
rect 20 32 22 36
<< ndiffusion >>
rect 6 8 10 12
rect 12 8 20 12
rect 22 8 26 12
<< pdiffusion >>
rect 6 32 10 36
rect 12 32 14 36
rect 18 32 20 36
rect 22 32 26 36
<< ndcontact >>
rect 2 8 6 12
rect 26 8 30 12
<< pdcontact >>
rect 2 32 6 36
rect 14 32 18 36
rect 26 32 30 36
<< psubstratepcontact >>
rect 2 0 6 4
<< nsubstratencontact >>
rect 2 40 6 44
rect 26 40 30 44
<< polysilicon >>
rect 10 36 12 38
rect 20 36 22 38
rect 10 24 12 32
rect 9 20 12 24
rect 10 12 12 20
rect 20 17 22 32
rect 19 13 22 17
rect 20 12 22 13
rect 10 6 12 8
rect 20 6 22 8
<< polycontact >>
rect 5 20 9 24
rect 15 13 19 17
<< metal1 >>
rect 0 40 2 44
rect 6 40 26 44
rect 30 40 32 44
rect 2 36 6 40
rect 26 36 30 40
rect 14 24 18 32
rect 14 20 30 24
rect 26 12 30 20
rect 2 4 6 8
rect 0 0 2 4
rect 6 0 32 4
<< labels >>
rlabel psubstratepcontact 4 2 4 2 1 VSS
rlabel nsubstratencontact 4 42 4 42 5 VDD
rlabel nsubstratencontact 28 42 28 42 5 VDD
rlabel polycontact 7 22 7 22 1 A
rlabel polycontact 17 15 17 15 1 B
rlabel metal1 28 22 28 22 1 Y
<< end >>
