magic
tech scmos
timestamp 1711474285
<< ntransistor >>
rect 4 -1 6 3
rect 26 -1 28 3
rect 44 -1 46 3
<< ptransistor >>
rect 4 39 6 43
rect 26 39 28 43
rect 44 39 46 43
<< ndiffusion >>
rect 2 -1 4 3
rect 6 -1 14 3
rect 18 -1 26 3
rect 28 -1 30 3
rect 42 -1 44 3
rect 46 -1 47 3
<< pdiffusion >>
rect 2 39 4 43
rect 6 39 26 43
rect 28 39 30 43
rect 42 39 44 43
rect 46 39 47 43
<< ndcontact >>
rect -2 -1 2 3
rect 14 -1 18 3
rect 30 -1 34 3
rect 38 -1 42 3
rect 47 -1 51 3
<< pdcontact >>
rect -2 39 2 43
rect 30 39 34 43
rect 38 39 42 43
rect 47 39 51 43
<< psubstratepcontact >>
rect -2 -9 2 -5
rect 30 -9 34 -5
rect 38 -9 42 -5
<< nsubstratencontact >>
rect -2 47 2 51
rect 38 47 42 51
<< polysilicon >>
rect 4 43 6 45
rect 26 43 28 45
rect 44 43 46 45
rect 4 11 6 39
rect 26 19 28 39
rect 24 15 28 19
rect 2 7 6 11
rect 4 3 6 7
rect 26 3 28 15
rect 44 11 46 39
rect 42 7 46 11
rect 44 3 46 7
rect 4 -4 6 -1
rect 26 -3 28 -1
rect 44 -3 46 -1
<< polycontact >>
rect 20 15 24 19
rect -2 7 2 11
rect 38 7 42 11
<< metal1 >>
rect -4 47 -2 51
rect 2 47 38 51
rect 42 47 53 51
rect -2 43 2 47
rect 38 43 42 47
rect 30 11 34 39
rect 14 7 38 11
rect 14 3 18 7
rect 47 3 51 39
rect -2 -5 2 -1
rect 30 -5 34 -1
rect 38 -5 42 -1
rect -4 -9 -2 -5
rect 2 -9 30 -5
rect 34 -9 38 -5
rect 42 -9 54 -5
<< labels >>
rlabel polycontact 0 9 0 9 1 A
rlabel polycontact 40 9 40 9 1 INV
rlabel metal1 49 10 49 10 1 Y
rlabel psubstratepcontact 0 -7 0 -7 1 VSS
rlabel psubstratepcontact 32 -7 32 -7 1 VSS
rlabel psubstratepcontact 40 -7 40 -7 1 VSS
rlabel polycontact 22 17 22 17 1 B
rlabel nsubstratencontact 0 49 0 49 4 VDD
<< end >>
