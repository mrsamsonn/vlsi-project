magic
tech scmos
timestamp 1707765594
<< nwell >>
rect -4 18 20 42
<< ntransistor >>
rect 7 8 9 12
<< ptransistor >>
rect 7 24 9 28
<< ndiffusion >>
rect 6 8 7 12
rect 9 8 10 12
<< pdiffusion >>
rect 6 24 7 28
rect 9 24 10 28
<< ndcontact >>
rect 2 8 6 12
rect 10 8 14 12
<< pdcontact >>
rect 2 24 6 28
rect 10 24 14 28
<< psubstratepcontact >>
rect 2 0 6 4
<< nsubstratencontact >>
rect 2 32 6 36
<< polysilicon >>
rect 7 28 9 30
rect 7 20 9 24
rect 6 16 9 20
rect 7 12 9 16
rect 7 6 9 8
<< polycontact >>
rect 2 16 6 20
<< metal1 >>
rect 0 32 2 36
rect 6 32 16 36
rect 2 28 6 32
rect 10 12 14 24
rect 2 4 6 8
rect 0 0 2 4
rect 6 0 16 4
<< labels >>
rlabel polycontact 4 17 4 17 1 A
rlabel metal1 12 17 12 17 1 Y
rlabel nsubstratencontact 4 34 4 34 1 VDD
rlabel psubstratepcontact 4 2 4 2 1 VSS
<< end >>
