magic
tech scmos
timestamp 1711520729
<< polycontact >>
rect 243 50 247 54
<< metal1 >>
rect 184 97 396 101
rect 92 89 260 93
rect 0 81 2 85
rect 182 81 186 85
rect 369 81 373 85
rect 274 53 286 57
rect 370 41 374 45
rect 423 37 427 73
rect 0 25 2 29
rect 183 25 187 29
rect 368 25 372 29
<< m2contact >>
rect 180 97 184 101
rect 396 97 400 101
rect 88 89 92 93
rect 260 89 264 93
rect 88 61 92 65
rect 180 61 184 65
rect 53 50 57 54
rect 74 50 78 54
rect 396 53 400 57
<< metal2 >>
rect 88 65 92 89
rect 180 65 184 97
rect 260 54 264 89
rect 396 57 400 97
use 2or  2or_0
timestamp 1711474285
transform 1 0 376 0 1 34
box -4 -9 54 51
use half-sub-2  half-sub-2_0
timestamp 1711519902
transform 1 0 186 0 1 0
box 0 0 184 85
use half-sub  half-sub_0
timestamp 1711519604
transform 1 0 0 0 1 0
box 0 0 184 85
<< labels >>
rlabel m2contact 55 52 55 52 1 B
rlabel m2contact 76 52 76 52 1 Bin
rlabel polycontact 245 52 245 52 1 A
rlabel metal1 425 54 425 54 7 Bout
rlabel metal1 280 55 280 55 1 Diff
rlabel metal1 1 83 1 83 3 VDD
rlabel metal1 1 27 1 27 3 VSS
<< end >>
