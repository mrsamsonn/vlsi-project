magic
tech scmos
timestamp 1710984200
<< ntransistor >>
rect 6 8 8 12
rect 20 8 22 12
rect 33 8 35 12
rect 54 8 56 12
<< ptransistor >>
rect 6 40 8 44
rect 20 40 22 44
rect 33 40 35 44
rect 54 40 56 44
<< ndiffusion >>
rect 4 8 6 12
rect 8 8 20 12
rect 22 8 24 12
rect 28 8 33 12
rect 35 8 54 12
rect 56 8 60 12
rect 64 8 68 12
<< pdiffusion >>
rect 4 40 6 44
rect 8 40 12 44
rect 16 40 20 44
rect 22 40 24 44
rect 28 40 33 44
rect 35 40 44 44
rect 48 40 54 44
rect 56 40 60 44
rect 64 40 68 44
<< ndcontact >>
rect 0 8 4 12
rect 24 8 28 12
rect 60 8 64 12
<< pdcontact >>
rect 0 40 4 44
rect 12 40 16 44
rect 24 40 28 44
rect 44 40 48 44
rect 60 40 64 44
<< psubstratepcontact >>
rect 24 0 28 4
<< nsubstratencontact >>
rect 12 56 16 60
<< polysilicon >>
rect 6 44 8 46
rect 20 44 22 46
rect 33 44 35 46
rect 54 44 56 46
rect 6 12 8 40
rect 20 12 22 40
rect 33 12 35 40
rect 54 12 56 40
rect 6 6 8 8
rect 20 6 22 8
rect 33 6 35 8
rect 54 6 56 8
<< polycontact >>
rect 2 25 6 29
rect 16 25 20 29
rect 29 25 33 29
rect 50 25 54 29
<< metal1 >>
rect -2 56 12 60
rect 16 56 70 60
rect 12 44 16 56
rect 24 48 64 52
rect 24 44 28 48
rect 60 44 64 48
rect 0 36 4 40
rect 24 36 28 40
rect 0 32 28 36
rect 44 36 48 40
rect 44 32 68 36
rect 60 20 64 32
rect 0 16 64 20
rect 0 12 4 16
rect 60 12 64 16
rect 24 4 28 8
rect -2 0 24 4
rect 28 0 70 4
<< labels >>
rlabel nsubstratencontact 14 58 14 58 5 VDD
rlabel psubstratepcontact 26 2 26 2 1 VSS
rlabel polycontact 4 27 4 27 3 A
rlabel polycontact 18 27 18 27 1 B
rlabel polycontact 31 27 31 27 1 B'
rlabel polycontact 52 27 52 27 1 A'
rlabel metal1 66 34 66 34 7 Y
<< end >>
